----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:05:29 11/22/2021 
-- Design Name: 
-- Module Name:    Sumador - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work_std_arith.all;

entity Sumador is
port (A, B : in std_logic_vector (0 to 1);
Z : out std_logic_vector (0 to 1));
end Sumador;

architecture Behavioral of Sumador is

begin


end Behavioral;

