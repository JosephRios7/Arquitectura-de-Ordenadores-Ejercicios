----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:04:41 11/22/2021 
-- Design Name: 
-- Module Name:    Bloque - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Bloque is
port (X: in std_logic_vector (1 downto 0);
A, B: in std_logic;
Z: out std_logic_vector (0 to 3));
end Bloque;

architecture Behavioral of Bloque is

begin


end Behavioral;

